1
0 0 0 0 0 r h 1 B 40 B 40 B 40 B
0 0 0 0 0 r h 12 B 53 B
0 0 0 0 0 r h 13 B 13 B 13 B 23 B 23 B
0 0 0 0 0 r h 32 B 45 B 45 B 45 B 32 B 32 B
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
4
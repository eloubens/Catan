3
4 1 1 3 0 r 16 19 36 h 15 T 27 H 36 B
0 3 2 4 2 r 11 17 h 10 T 50 T 38 T
3 2 2 2 3 r 43 0 1 h 29 H 34 H
3 2 0 3 0 r h 22 H
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
5
3
3 3 3 3 3 r 9 h 1 B 3 B
4 4 4 4 4 r 44 h 10 B 15 B 19 T
4 3 6 2 4 r 5 h 33 B 
1 3 5 7 9 r 33 70 h 19 H
0 3 1 10 3 5 1 4 5 7 3 10 5 7 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 5 7 4 6 2 9 2 9
17
0
0 0 0 0 0 r h 1 B
0 0 0 0 0 r h 3 B 3 B
0 0 0 0 0 r h
0 0 0 0 0 r h
3 5 2 11 3 12 1 9 2 4 2 11 1 8 1 2 3 4 0 3 0 6 4 8 4 9 2 3 4 7 0 6 1 5 5 10 0 10
17
1
0 0 0 0 1 r h 1 B 14 B
0 0 0 0 1 r h 3 B 12 B
0 0 0 0 0 r h 5 B 11 B
0 0 0 0 1 r h 7 B 9 B
4 10 0 3 1 8 2 6 1 6 2 7 5 8 3 9 1 9 4 11 0 5 1 3 2 12 2 5 3 10 0 2 4 4 3 4 0 11
6
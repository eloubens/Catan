0
0 0 0 0 0 r h 0 B
0 0 0 0 0 r h 4 B
0 0 0 0 0 r h
0 0 0 0 0 r h
0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0
0
0
0 0 0 0 0 r h 1 B
0 0 0 0 0 r h 3 B 3 B
0 0 0 0 0 r h 5 B
0 0 0 0 0 r h
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9
4